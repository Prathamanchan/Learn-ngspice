v1 1 0 150v
R1 1 2 20
R2 2 0 10
R3 2 3 15
V2 3 0 100V

.op
.end
