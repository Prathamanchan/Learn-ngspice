Ex3

G1 1 3 1 0 0.1  ;Voltage dependent current source
*G nodes of CS nodes of Dependent voltage - Dependence scale
R1 1 0 10
I1 0 2 10A
R2 1 2 5
R3 2 3 10
R4 3 0 5

.op
.end
