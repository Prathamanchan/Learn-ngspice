I-VCharacteristics of CD4007 
*Including the CD4007 model file
.include cd4007.txt
*Fixing gate bias at 3.5V
vgg 1 0 dc 3.5v
rg 1 2 680
*Specifying NMOS in this manner-
*name drain gate source body modelname
m1 3 2 0 0 MbreakND
rd 3 4 100
*DC analysis to sweep vds from 0 to 5
.dc vdd 0 5 0.01
.control
run
plot vid#branch vs v(3)
.endc
.end
